[aimspice]
[description]
3320
Untitled circuit* This is a parametrized testbench for your pixel circuit array

* You should at least test your circuit with:
*	- current of 50 pA and exposure time 30 ms
*	- current of 750 pA and exposure time 2 ms

* Instructions
* Connect EXPOSE, ERASE, NRE_R1 and NRE_R2 at the right place
* Run a transient simulation with length 60 ms
* Make sure outputs of pixel circuits to ADC are called OUT1 and OUT2
* Make plots of output voltages to ADC (here called OUT1 and OUT2)
* The voltage across internal capacitor (any pixel) is also of interest (here called OUT_SAMPLED1)
* You should also plot the control signals EXPOSE, NRE_R1, NRE_R2 and ERASE

.include PhotoDiode.cir
.include p18_model_card.inc
.include p18_cmos_models_tt.inc



.param Ipd_1 = 50p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 30m ! Exposusre time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency 
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param NRE_R2_DLY = {4*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R2 signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

VDD 1 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R1 NRE_R1 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R2 NRE_R2 0 dc 0  pulse(VDD 0 NRE_R2_DLY TRF TRF CLK_PERIOD PERIOD)

.subckt PixelSegment VDD VSS EXPOSE OUT
	xPD0 VDD OUT PhotoDiode Ipd=750p

	*DRAIN GATE  SOURCE BULK
	MN1 N1 EXPOSE OUT VSS NMOS L=2U W=2U
	
	!MN2 OUT ERASE VSS VSS NMOS L =0.7U W=3U
	
	C1 OUT VSS 1u	
	!R0 OUT VSS 1k

.ends
		******************
		***DEFINE PIXEL***
		******************
 
.subckt Pixel VDD VSS EXPOSE ERASE NRE OUT
	xPD1 VDD N1 PhotoDiode Ipd=750p

	*DRAIN GATE  SOURCE BULK
	M1 N1 EXPOSE N2 VSS NMOS L=0.36U W=5.04U
	
	M2 N2 ERASE VSS VSS NMOS L =1.08U W=1.08U
	
	C1 N2 VSS 2p	

	M3 VSS N2 N3 VDD PMOS L =0.36U W=5.04U
	M4 N3 NRE OUT VDD PMOS L =1.08U W=1.08U
	!R0 OUT VDD 10M
.ends 

		************************
		***DEFINE PIXEL ARRAY***
		************************

.subckt PixelArray VDD VSS EXPOSE ERASE NRE_R1 NRE_R2 OUT1 OUT2
	
	**PIXEL**
	xPixel1_1 VDD VSS EXPOSE ERASE NRE_R1 OUT1 Pixel
	xPixel1_2 VDD VSS EXPOSE ERASE NRE_R1 OUT2 Pixel
	xPixel2_1 VDD VSS EXPOSE ERASE NRE_R2 OUT1 Pixel
	xPixel2_2 VDD VSS EXPOSE ERASE NRE_R2 OUT2 Pixel

	**LOAD**
	MC1 OUT1 OUT1 VDD VDD PMOS L =1.0U W=1.67U
	MC2 OUT2 OUT2 VDD VDD PMOS L =1.0U W=1.67U

	**CAPACITORS**
	CC1 OUT1 VSS 3p
	CC2 OUT1 VSS 3p

.ends

xmy_pixelArray 1 0 EXPOSE ERASE NRE_R1 NRE_R2 OUT1 OUT2 PixelArray


!xmy_pixel 1 0 EXPOSE ERASE NRE_R1 OUT Pixel
!.plot V(OUT)


.plot V(EXPOSE) V(ERASE) V(NRE_R1) V(OUT1)
!.plot V(OUT1) V(OUT2) ! signals going to ADC
!.plot V(EXPOSE) V(NRE_R1) V(NRE_R2) V(ERASE)
!.plot V(OUT_SAMPLED1)
[dc]
1
V1
1
3
0.1
[tran]
0.1m
60m
X
X
0
[ana]
4 0
[end]
